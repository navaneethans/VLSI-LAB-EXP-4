6(iii): D FLIP FLOP 
module dff( clk,d,q); 
input clk,d; 
output reg q; 



endmodule