6(iv):T FLIPFLOP 
module tff(t,clk,q); 
input t,clk; 
output reg q=1; 



endmodule