module sr( s,r,clk,q);
 input s,r,clk; 
output reg q=0; 




endmodule





