6(ii): JK FLIP FLOP 
module jk( j,k,clk,q); 
input j,k,clk; 
output reg q=0; 



endmodule